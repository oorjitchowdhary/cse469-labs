// 64 bit program counter
